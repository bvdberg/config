library ieee;
use ieee.std_logic_1164.all;

entity AbcTb is
end entity;

architecture sim of AcbTb is

begin

    process is
    begin

        wait for 10 ns;

    end process;

end architecture;

